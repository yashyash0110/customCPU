`define ADD   = 5'b00000
`define SUB   = 5'b00001
`define MUL   = 5'b00010
`define DIV   = 5'b00011
`define INC   = 5'b00100
`define DEC   = 5'b00101
`define AND   = 5'b00110
`define OR    = 5'b00111
`define XOR   = 5'b01000
`define NOT   = 5'b01001
`define JMP   = 5'b01010
`define BEQ   = 5'b01011
`define BNE   = 5'b01100
`define CALL  = 5'b01101
`define RET   = 5'b01110
`define LD    = 5'b01111
`define ST    = 5'b10000
`define FFT   = 5'b10001
`define ENC   = 5'b10010
`define DEC2  = 5'b10011
